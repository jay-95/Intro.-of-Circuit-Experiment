module Segment_str (s,A,B);
  
endmodule