library verilog;
use verilog.vl_types.all;
entity tb_Encoder_4X2 is
end tb_Encoder_4X2;
