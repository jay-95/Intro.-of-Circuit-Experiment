`timescale 1ns/10ps
module tb_Segment;
  reg B,A;
  wire [0:6] sdout;
  wire [0:3] D;
  
  BCD_to_7_Segment_Decoder u1(sdout,D);
  Decoder_2X4 u2(D,A,B);
    
  initial
  begin
    B = 1'b0;
    A = 1'b0;
    
    #10 A = 1'b1;
    
    #10 B = 1'b1;
        A = 1'b0;
    
    #10 A = 1'b1`timescale 1ns/10ps
module tb_Segment;
  reg B,A;
  wire [0:6] sdout;
  wire [0:3] D;
  
  BCD_to_7_Segment_Decoder u1(sdout,D);
  Decoder_2X4 u2(D,A,B);
    
  initial
  begin
    B = 1'b0;
    A = 1'b0;
    
    #10 A = 1'b1;
    
    #10 B = 1'b1;
        A = 1'b0;
    
    #10 A = 1'b1;
    
    #10 $stop;
  end
endmodule;
    
    #10 $stop;
  end
endmodule