library verilog;
use verilog.vl_types.all;
entity tb_ripple is
end tb_ripple;
