library verilog;
use verilog.vl_types.all;
entity tb_Decoder_2X4 is
end tb_Decoder_2X4;
