library verilog;
use verilog.vl_types.all;
entity tb_Segment is
end tb_Segment;
